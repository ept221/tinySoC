module test_tb();

    reg clk = 0;

endmodule